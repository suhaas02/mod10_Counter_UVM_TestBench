package counter_test_pkg;  

	import uvm_pkg::*;
	`include "uvm_macros.svh"
   	//`include the files 
	`include "transaction.sv"
	`include "count_config.sv"
 	`include "driver.sv"
 	`include "monitor.sv"
	`include "sequencer.sv"
	`include "agent.sv" 
 	`include "scoreboard.sv"
 	`include "environment.sv"
	`include "sequence.sv"
 	`include "test.sv" 
endpackage
	
